`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   00:08:05 09/28/2020
// Design Name:   fba
// Module Name:   D:/College/CS/F215/Exp_6_2019A7PS0097H/four_adder.v
// Project Name:  Exp_6_2019A7PS0097H
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: fba
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module four_adder;

	// Inputs
	reg [3:0] A;
	reg [3:0] B;

	// Outputs
	wire [3:0] Sum;
	wire Carry;

	// Instantiate the Unit Under Test (UUT)
	fba uut (
		.A(A), 
		.B(B), 
		.Sum(Sum), 
		.Carry(Carry)
	);

	initial begin

		A = 0 ;
		B = 0 ;
		#1 ;

		A = 0 ;
		B = 1 ;
		#1 ;

		A = 0 ;
		B = 2 ;
		#1 ;

		A = 0 ;
		B = 3 ;
		#1 ;

		A = 0 ;
		B = 4 ;
		#1 ;

		A = 0 ;
		B = 5 ;
		#1 ;

		A = 0 ;
		B = 6 ;
		#1 ;

		A = 0 ;
		B = 7 ;
		#1 ;

		A = 0 ;
		B = 8 ;
		#1 ;

		A = 0 ;
		B = 9 ;
		#1 ;

		A = 0 ;
		B = 10 ;
		#1 ;

		A = 0 ;
		B = 11 ;
		#1 ;

		A = 0 ;
		B = 12 ;
		#1 ;

		A = 0 ;
		B = 13 ;
		#1 ;

		A = 0 ;
		B = 14 ;
		#1 ;

		A = 0 ;
		B = 15 ;
		#1 ;


		A = 1 ;
		B = 0 ;
		#1 ;

		A = 1 ;
		B = 1 ;
		#1 ;

		A = 1 ;
		B = 2 ;
		#1 ;

		A = 1 ;
		B = 3 ;
		#1 ;

		A = 1 ;
		B = 4 ;
		#1 ;

		A = 1 ;
		B = 5 ;
		#1 ;

		A = 1 ;
		B = 6 ;
		#1 ;

		A = 1 ;
		B = 7 ;
		#1 ;

		A = 1 ;
		B = 8 ;
		#1 ;

		A = 1 ;
		B = 9 ;
		#1 ;

		A = 1 ;
		B = 10 ;
		#1 ;

		A = 1 ;
		B = 11 ;
		#1 ;

		A = 1 ;
		B = 12 ;
		#1 ;

		A = 1 ;
		B = 13 ;
		#1 ;

		A = 1 ;
		B = 14 ;
		#1 ;

		A = 1 ;
		B = 15 ;
		#1 ;


		A = 2 ;
		B = 0 ;
		#1 ;

		A = 2 ;
		B = 1 ;
		#1 ;

		A = 2 ;
		B = 2 ;
		#1 ;

		A = 2 ;
		B = 3 ;
		#1 ;

		A = 2 ;
		B = 4 ;
		#1 ;

		A = 2 ;
		B = 5 ;
		#1 ;

		A = 2 ;
		B = 6 ;
		#1 ;

		A = 2 ;
		B = 7 ;
		#1 ;

		A = 2 ;
		B = 8 ;
		#1 ;

		A = 2 ;
		B = 9 ;
		#1 ;

		A = 2 ;
		B = 10 ;
		#1 ;

		A = 2 ;
		B = 11 ;
		#1 ;

		A = 2 ;
		B = 12 ;
		#1 ;

		A = 2 ;
		B = 13 ;
		#1 ;

		A = 2 ;
		B = 14 ;
		#1 ;

		A = 2 ;
		B = 15 ;
		#1 ;


		A = 3 ;
		B = 0 ;
		#1 ;

		A = 3 ;
		B = 1 ;
		#1 ;

		A = 3 ;
		B = 2 ;
		#1 ;

		A = 3 ;
		B = 3 ;
		#1 ;

		A = 3 ;
		B = 4 ;
		#1 ;

		A = 3 ;
		B = 5 ;
		#1 ;

		A = 3 ;
		B = 6 ;
		#1 ;

		A = 3 ;
		B = 7 ;
		#1 ;

		A = 3 ;
		B = 8 ;
		#1 ;

		A = 3 ;
		B = 9 ;
		#1 ;

		A = 3 ;
		B = 10 ;
		#1 ;

		A = 3 ;
		B = 11 ;
		#1 ;

		A = 3 ;
		B = 12 ;
		#1 ;

		A = 3 ;
		B = 13 ;
		#1 ;

		A = 3 ;
		B = 14 ;
		#1 ;

		A = 3 ;
		B = 15 ;
		#1 ;


		A = 4 ;
		B = 0 ;
		#1 ;

		A = 4 ;
		B = 1 ;
		#1 ;

		A = 4 ;
		B = 2 ;
		#1 ;

		A = 4 ;
		B = 3 ;
		#1 ;

		A = 4 ;
		B = 4 ;
		#1 ;

		A = 4 ;
		B = 5 ;
		#1 ;

		A = 4 ;
		B = 6 ;
		#1 ;

		A = 4 ;
		B = 7 ;
		#1 ;

		A = 4 ;
		B = 8 ;
		#1 ;

		A = 4 ;
		B = 9 ;
		#1 ;

		A = 4 ;
		B = 10 ;
		#1 ;

		A = 4 ;
		B = 11 ;
		#1 ;

		A = 4 ;
		B = 12 ;
		#1 ;

		A = 4 ;
		B = 13 ;
		#1 ;

		A = 4 ;
		B = 14 ;
		#1 ;

		A = 4 ;
		B = 15 ;
		#1 ;


		A = 5 ;
		B = 0 ;
		#1 ;

		A = 5 ;
		B = 1 ;
		#1 ;

		A = 5 ;
		B = 2 ;
		#1 ;

		A = 5 ;
		B = 3 ;
		#1 ;

		A = 5 ;
		B = 4 ;
		#1 ;

		A = 5 ;
		B = 5 ;
		#1 ;

		A = 5 ;
		B = 6 ;
		#1 ;

		A = 5 ;
		B = 7 ;
		#1 ;

		A = 5 ;
		B = 8 ;
		#1 ;

		A = 5 ;
		B = 9 ;
		#1 ;

		A = 5 ;
		B = 10 ;
		#1 ;

		A = 5 ;
		B = 11 ;
		#1 ;

		A = 5 ;
		B = 12 ;
		#1 ;

		A = 5 ;
		B = 13 ;
		#1 ;

		A = 5 ;
		B = 14 ;
		#1 ;

		A = 5 ;
		B = 15 ;
		#1 ;


		A = 6 ;
		B = 0 ;
		#1 ;

		A = 6 ;
		B = 1 ;
		#1 ;

		A = 6 ;
		B = 2 ;
		#1 ;

		A = 6 ;
		B = 3 ;
		#1 ;

		A = 6 ;
		B = 4 ;
		#1 ;

		A = 6 ;
		B = 5 ;
		#1 ;

		A = 6 ;
		B = 6 ;
		#1 ;

		A = 6 ;
		B = 7 ;
		#1 ;

		A = 6 ;
		B = 8 ;
		#1 ;

		A = 6 ;
		B = 9 ;
		#1 ;

		A = 6 ;
		B = 10 ;
		#1 ;

		A = 6 ;
		B = 11 ;
		#1 ;

		A = 6 ;
		B = 12 ;
		#1 ;

		A = 6 ;
		B = 13 ;
		#1 ;

		A = 6 ;
		B = 14 ;
		#1 ;

		A = 6 ;
		B = 15 ;
		#1 ;


		A = 7 ;
		B = 0 ;
		#1 ;

		A = 7 ;
		B = 1 ;
		#1 ;

		A = 7 ;
		B = 2 ;
		#1 ;

		A = 7 ;
		B = 3 ;
		#1 ;

		A = 7 ;
		B = 4 ;
		#1 ;

		A = 7 ;
		B = 5 ;
		#1 ;

		A = 7 ;
		B = 6 ;
		#1 ;

		A = 7 ;
		B = 7 ;
		#1 ;

		A = 7 ;
		B = 8 ;
		#1 ;

		A = 7 ;
		B = 9 ;
		#1 ;

		A = 7 ;
		B = 10 ;
		#1 ;

		A = 7 ;
		B = 11 ;
		#1 ;

		A = 7 ;
		B = 12 ;
		#1 ;

		A = 7 ;
		B = 13 ;
		#1 ;

		A = 7 ;
		B = 14 ;
		#1 ;

		A = 7 ;
		B = 15 ;
		#1 ;


		A = 8 ;
		B = 0 ;
		#1 ;

		A = 8 ;
		B = 1 ;
		#1 ;

		A = 8 ;
		B = 2 ;
		#1 ;

		A = 8 ;
		B = 3 ;
		#1 ;

		A = 8 ;
		B = 4 ;
		#1 ;

		A = 8 ;
		B = 5 ;
		#1 ;

		A = 8 ;
		B = 6 ;
		#1 ;

		A = 8 ;
		B = 7 ;
		#1 ;

		A = 8 ;
		B = 8 ;
		#1 ;

		A = 8 ;
		B = 9 ;
		#1 ;

		A = 8 ;
		B = 10 ;
		#1 ;

		A = 8 ;
		B = 11 ;
		#1 ;

		A = 8 ;
		B = 12 ;
		#1 ;

		A = 8 ;
		B = 13 ;
		#1 ;

		A = 8 ;
		B = 14 ;
		#1 ;

		A = 8 ;
		B = 15 ;
		#1 ;


		A = 9 ;
		B = 0 ;
		#1 ;

		A = 9 ;
		B = 1 ;
		#1 ;

		A = 9 ;
		B = 2 ;
		#1 ;

		A = 9 ;
		B = 3 ;
		#1 ;

		A = 9 ;
		B = 4 ;
		#1 ;

		A = 9 ;
		B = 5 ;
		#1 ;

		A = 9 ;
		B = 6 ;
		#1 ;

		A = 9 ;
		B = 7 ;
		#1 ;

		A = 9 ;
		B = 8 ;
		#1 ;

		A = 9 ;
		B = 9 ;
		#1 ;

		A = 9 ;
		B = 10 ;
		#1 ;

		A = 9 ;
		B = 11 ;
		#1 ;

		A = 9 ;
		B = 12 ;
		#1 ;

		A = 9 ;
		B = 13 ;
		#1 ;

		A = 9 ;
		B = 14 ;
		#1 ;

		A = 9 ;
		B = 15 ;
		#1 ;


		A = 10 ;
		B = 0 ;
		#1 ;

		A = 10 ;
		B = 1 ;
		#1 ;

		A = 10 ;
		B = 2 ;
		#1 ;

		A = 10 ;
		B = 3 ;
		#1 ;

		A = 10 ;
		B = 4 ;
		#1 ;

		A = 10 ;
		B = 5 ;
		#1 ;

		A = 10 ;
		B = 6 ;
		#1 ;

		A = 10 ;
		B = 7 ;
		#1 ;

		A = 10 ;
		B = 8 ;
		#1 ;

		A = 10 ;
		B = 9 ;
		#1 ;

		A = 10 ;
		B = 10 ;
		#1 ;

		A = 10 ;
		B = 11 ;
		#1 ;

		A = 10 ;
		B = 12 ;
		#1 ;

		A = 10 ;
		B = 13 ;
		#1 ;

		A = 10 ;
		B = 14 ;
		#1 ;

		A = 10 ;
		B = 15 ;
		#1 ;


		A = 11 ;
		B = 0 ;
		#1 ;

		A = 11 ;
		B = 1 ;
		#1 ;

		A = 11 ;
		B = 2 ;
		#1 ;

		A = 11 ;
		B = 3 ;
		#1 ;

		A = 11 ;
		B = 4 ;
		#1 ;

		A = 11 ;
		B = 5 ;
		#1 ;

		A = 11 ;
		B = 6 ;
		#1 ;

		A = 11 ;
		B = 7 ;
		#1 ;

		A = 11 ;
		B = 8 ;
		#1 ;

		A = 11 ;
		B = 9 ;
		#1 ;

		A = 11 ;
		B = 10 ;
		#1 ;

		A = 11 ;
		B = 11 ;
		#1 ;

		A = 11 ;
		B = 12 ;
		#1 ;

		A = 11 ;
		B = 13 ;
		#1 ;

		A = 11 ;
		B = 14 ;
		#1 ;

		A = 11 ;
		B = 15 ;
		#1 ;


		A = 12 ;
		B = 0 ;
		#1 ;

		A = 12 ;
		B = 1 ;
		#1 ;

		A = 12 ;
		B = 2 ;
		#1 ;

		A = 12 ;
		B = 3 ;
		#1 ;

		A = 12 ;
		B = 4 ;
		#1 ;

		A = 12 ;
		B = 5 ;
		#1 ;

		A = 12 ;
		B = 6 ;
		#1 ;

		A = 12 ;
		B = 7 ;
		#1 ;

		A = 12 ;
		B = 8 ;
		#1 ;

		A = 12 ;
		B = 9 ;
		#1 ;

		A = 12 ;
		B = 10 ;
		#1 ;

		A = 12 ;
		B = 11 ;
		#1 ;

		A = 12 ;
		B = 12 ;
		#1 ;

		A = 12 ;
		B = 13 ;
		#1 ;

		A = 12 ;
		B = 14 ;
		#1 ;

		A = 12 ;
		B = 15 ;
		#1 ;


		A = 13 ;
		B = 0 ;
		#1 ;

		A = 13 ;
		B = 1 ;
		#1 ;

		A = 13 ;
		B = 2 ;
		#1 ;

		A = 13 ;
		B = 3 ;
		#1 ;

		A = 13 ;
		B = 4 ;
		#1 ;

		A = 13 ;
		B = 5 ;
		#1 ;

		A = 13 ;
		B = 6 ;
		#1 ;

		A = 13 ;
		B = 7 ;
		#1 ;

		A = 13 ;
		B = 8 ;
		#1 ;

		A = 13 ;
		B = 9 ;
		#1 ;

		A = 13 ;
		B = 10 ;
		#1 ;

		A = 13 ;
		B = 11 ;
		#1 ;

		A = 13 ;
		B = 12 ;
		#1 ;

		A = 13 ;
		B = 13 ;
		#1 ;

		A = 13 ;
		B = 14 ;
		#1 ;

		A = 13 ;
		B = 15 ;
		#1 ;


		A = 14 ;
		B = 0 ;
		#1 ;

		A = 14 ;
		B = 1 ;
		#1 ;

		A = 14 ;
		B = 2 ;
		#1 ;

		A = 14 ;
		B = 3 ;
		#1 ;

		A = 14 ;
		B = 4 ;
		#1 ;

		A = 14 ;
		B = 5 ;
		#1 ;

		A = 14 ;
		B = 6 ;
		#1 ;

		A = 14 ;
		B = 7 ;
		#1 ;

		A = 14 ;
		B = 8 ;
		#1 ;

		A = 14 ;
		B = 9 ;
		#1 ;

		A = 14 ;
		B = 10 ;
		#1 ;

		A = 14 ;
		B = 11 ;
		#1 ;

		A = 14 ;
		B = 12 ;
		#1 ;

		A = 14 ;
		B = 13 ;
		#1 ;

		A = 14 ;
		B = 14 ;
		#1 ;

		A = 14 ;
		B = 15 ;
		#1 ;


		A = 15 ;
		B = 0 ;
		#1 ;

		A = 15 ;
		B = 1 ;
		#1 ;

		A = 15 ;
		B = 2 ;
		#1 ;

		A = 15 ;
		B = 3 ;
		#1 ;

		A = 15 ;
		B = 4 ;
		#1 ;

		A = 15 ;
		B = 5 ;
		#1 ;

		A = 15 ;
		B = 6 ;
		#1 ;

		A = 15 ;
		B = 7 ;
		#1 ;

		A = 15 ;
		B = 8 ;
		#1 ;

		A = 15 ;
		B = 9 ;
		#1 ;

		A = 15 ;
		B = 10 ;
		#1 ;

		A = 15 ;
		B = 11 ;
		#1 ;

		A = 15 ;
		B = 12 ;
		#1 ;

		A = 15 ;
		B = 13 ;
		#1 ;

		A = 15 ;
		B = 14 ;
		#1 ;

		A = 15 ;
		B = 15 ;
		#1 ;
		
		$finish ;

	end
      
endmodule

