`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   08:46:12 10/27/2020
// Design Name:   Mux
// Module Name:   D:/College/CS/F215/Exp_9_2019A7PS0097H/muxtest.v
// Project Name:  Exp_9_2019A7PS0097H
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Mux
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module muxtest;

	// Inputs
	reg [7:0] I;
	reg [2:0] S;

	// Outputs
	wire Y;

	// Instantiate the Unit Under Test (UUT)
	Mux uut (
		.I(I), 
		.S(S), 
		.Y(Y)
	);

	initial begin
		
		I = 0000000 ;
		S = 000 ;
		$10 ;

		I = 0000000 ;
		S = 001 ;
		$10 ;

		I = 0000000 ;
		S = 010 ;
		$10 ;

		I = 0000000 ;
		S = 011 ;
		$10 ;

		I = 0000000 ;
		S = 100 ;
		$10 ;

		I = 0000000 ;
		S = 101 ;
		$10 ;

		I = 0000000 ;
		S = 110 ;
		$10 ;

		I = 0000000 ;
		S = 111 ;
		$10 ;

		I = 0000001 ;
		S = 000 ;
		$10 ;

		I = 0000001 ;
		S = 001 ;
		$10 ;

		I = 0000001 ;
		S = 010 ;
		$10 ;

		I = 0000001 ;
		S = 011 ;
		$10 ;

		I = 0000001 ;
		S = 100 ;
		$10 ;

		I = 0000001 ;
		S = 101 ;
		$10 ;

		I = 0000001 ;
		S = 110 ;
		$10 ;

		I = 0000001 ;
		S = 111 ;
		$10 ;

		I = 0000010 ;
		S = 000 ;
		$10 ;

		I = 0000010 ;
		S = 001 ;
		$10 ;

		I = 0000010 ;
		S = 010 ;
		$10 ;

		I = 0000010 ;
		S = 011 ;
		$10 ;

		I = 0000010 ;
		S = 100 ;
		$10 ;

		I = 0000010 ;
		S = 101 ;
		$10 ;

		I = 0000010 ;
		S = 110 ;
		$10 ;

		I = 0000010 ;
		S = 111 ;
		$10 ;

		I = 0000100 ;
		S = 000 ;
		$10 ;

		I = 0000100 ;
		S = 001 ;
		$10 ;

		I = 0000100 ;
		S = 010 ;
		$10 ;

		I = 0000100 ;
		S = 011 ;
		$10 ;

		I = 0000100 ;
		S = 100 ;
		$10 ;

		I = 0000100 ;
		S = 101 ;
		$10 ;

		I = 0000100 ;
		S = 110 ;
		$10 ;

		I = 0000100 ;
		S = 111 ;
		$10 ;

		I = 0001000 ;
		S = 000 ;
		$10 ;

		I = 0001000 ;
		S = 001 ;
		$10 ;

		I = 0001000 ;
		S = 010 ;
		$10 ;

		I = 0001000 ;
		S = 011 ;
		$10 ;

		I = 0001000 ;
		S = 100 ;
		$10 ;

		I = 0001000 ;
		S = 101 ;
		$10 ;

		I = 0001000 ;
		S = 110 ;
		$10 ;

		I = 0001000 ;
		S = 111 ;
		$10 ;

		I = 0010000 ;
		S = 000 ;
		$10 ;

		I = 0010000 ;
		S = 001 ;
		$10 ;

		I = 0010000 ;
		S = 010 ;
		$10 ;

		I = 0010000 ;
		S = 011 ;
		$10 ;

		I = 0010000 ;
		S = 100 ;
		$10 ;

		I = 0010000 ;
		S = 101 ;
		$10 ;

		I = 0010000 ;
		S = 110 ;
		$10 ;

		I = 0010000 ;
		S = 111 ;
		$10 ;

		I = 0100000 ;
		S = 000 ;
		$10 ;

		I = 0100000 ;
		S = 001 ;
		$10 ;

		I = 0100000 ;
		S = 010 ;
		$10 ;

		I = 0100000 ;
		S = 011 ;
		$10 ;

		I = 0100000 ;
		S = 100 ;
		$10 ;

		I = 0100000 ;
		S = 101 ;
		$10 ;

		I = 0100000 ;
		S = 110 ;
		$10 ;

		I = 0100000 ;
		S = 111 ;
		$10 ;

		I = 1000000 ;
		S = 000 ;
		$10 ;

		I = 1000000 ;
		S = 001 ;
		$10 ;

		I = 1000000 ;
		S = 010 ;
		$10 ;

		I = 1000000 ;
		S = 011 ;
		$10 ;

		I = 1000000 ;
		S = 100 ;
		$10 ;

		I = 1000000 ;
		S = 101 ;
		$10 ;

		I = 1000000 ;
		S = 110 ;
		$10 ;

		I = 1000000 ;
		S = 111 ;
		$10 ;
		
		$finish ;

			end
      
endmodule

